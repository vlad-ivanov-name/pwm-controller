module clock_synchronizer (
	input wire in_clk_i,
	input wire out_clk_i,
	
	input wire data_i,
	output reg data_o
);

endmodule